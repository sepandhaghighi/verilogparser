// Verilog
// c17
// Ninputs 5
// Noutputs 2
// NtotalGates 6
// NAND2 6

module c17 (N1,N2,N3);

input N1,N2;

output N3;


or NAND2_1 (N3, N1, N2);


endmodule
