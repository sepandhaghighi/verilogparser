module c17 (N1,N2,N3);

input N1,N2;

output N3;


xor NAND2_1 (N3,N1,N2);

endmodule